//0613246
//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;

//Sign extended

always @ (data_i) begin

	data_o[16-1:0] = data_i;

	if(data_o[15]==1)
		data_o[32-1:16]=16'd65535;
	else
		data_o[32-1:16]=16'd0;
end
          
endmodule      
     